

module top(

    );
endmodule
