`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/30/2025 12:35:41 PM
// Design Name: 
// Module Name: alu
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module alu (
    input [31:0] a, b,                // Operands (32-bit by default)
    input [2:0] ALUControl,           // Selects ALU operation
    output reg [31:0] Result,         // Result of ALU operation
    output Zero,                      // 1 if Result is zero
    input funct7bit6,                 // Used to distinguish SRL vs SRA
    input funct3_bit                  // Used to distinguish SLT vs SLTU
);


always @(*) begin
    case(ALUControl)
        3'b000: Result = a + b; //add
        3'b001: Result = a - b; //sub
        3'b010: Result = a & b; //and
        3'b011: Result = a | b; //or
        3'b100: Result = a << b[4:0]; //sll
        
        
        
        3'b101: case (funct3_bit)

            1'b0:begin//slt
                if(a[31]!= b[31]) Result = a[31] ?1:0; 
                else Result = (a < b) ? 1:0;
            end 
            1'b1: Result <= (a < {20'b0, b[11:0]}) ? 1 : 0; //sltu
                endcase
                
                
        3'b110: begin
            if(funct7bit6) Result = a >> b[4:0]; //srl
            else Result = a >>> b[4:0]; //sra
        end
        
        
        
        3'b111: Result = a ^ b; //xor
        default: Result = 32'b0;
        endcase
end

assign Zero = (Result == 0)?1:0;

endmodule

/*
module alu(a,b,ALUcontrol,result,zero,negative,overflow,carry);
    input [31:0] a,b;       //two 32-bit inputs (operands)
    input [2:0] ALUcontrol; //control signals to determine the operation required 
                            //8 operations possible
    output [31:0] result;   //32-bit result
    
    output zero,negative,overflow,carry;
    
    //considering there will be a presence of internal wires
    //datapath declaration
    wire [31:0] a_and_b;
    wire [31:0] a_or_b;
    wire [31:0] not_b;
    
    wire [31:0] mux_res;
    
    wire [31:0] final_mux_res;
    
    wire [32:0] full_sum;
    wire [31:0] sum;
    wire cout;
    
    wire [31:0] slt; //set less than operation
    
    wire add_overflow;
    wire sub_overflow;
    
    
    //main logic
    
    //AND operation
    assign a_and_b = a & b;
    
    //OR operation
    assign a_or_b = a | b;
    
    //NOT operation
    assign not_b = ~b; 
    
    //mux operation 
    assign mux_res = (ALUcontrol[0] == 1'b0) ? b : not_b;
    //ALUcontrol is a 3 bit register, so one bit (0th) is taken from it to for bit extraction
    
    assign full_sum = a + mux_res + ALUcontrol[0]; //ALUControl[0]=0, then sum
                                                        //ALUControl[0]=1, them subtraction (2's complement)
                                                        
    assign sum = full_sum[31:0];
    assign cout = full_sum[32];                         //cout = 1, if addition results in 33 bit
                                                        //cout = 0, if addition results in 32 bit
    
   
    //Zero extension
    assign slt = {31'b0000000000000000000000000000000,sum[31]};    
    
    //final alu result logic
    assign final_mux_res = (ALUcontrol[2:0] == 3'b000) ? sum : //sum of a + b
                           (ALUcontrol[2:0] == 3'b001) ? sum : //sum of a + (-b) (subtraction)
                           (ALUcontrol[2:0] == 3'b010) ? a_and_b : 
                           (ALUcontrol[2:0] == 3'b011) ? a_or_b :
                           (ALUcontrol[2:0] == 3'b101) ? slt : 32'h00000000;
                         
    assign result = final_mux_res; //final result generation
    
    
    //flags 
    assign zero = (result == 32'b0);   //~result & ~result  
    assign negative = result[31]; //1:-ve, 0:+ve
    assign carry = (ALUcontrol == 3'b000) ? cout : 1'b0; //carry generated by the result
    
    
    // For a + b overflow
    assign add_overflow = (~a[31] & ~b[31] & sum[31]) | (a[31] & b[31] & ~sum[31]);
    
    // For a - b overflow
    // Subtraction is a + (-b), so signs are different
    assign sub_overflow = (~a[31] & b[31] & sum[31]) | (a[31] & ~b[31] & ~sum[31]);
    
    // Use ALU control to pick the correct one
    assign overflow = (ALUcontrol == 3'b000) ? add_overflow :
                      (ALUcontrol == 3'b001) ? sub_overflow : 1'b0;
                      
    
endmodule
*/
